library ieee;
use ieee.std 


enitity full
